module dut(input reg a,
	input reg b,
	output wire y
);
assign y=a^b;
endmodule
